module top_module (
    input clk,
    input [7:0] in,
    output reg [7:0]pedge
);
    wire [7:0] last;
    always@(posedge clk) 
        begin
            pedge <= ~last&in; 
            last <= in;
        end
endmodule
